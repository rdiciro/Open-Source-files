* SPICE3 file created from layout_test1.ext - technology: sky130A

X0 XM2/vdd XM2/vin XM2/vout XM2/vdd sky130_fd_pr__pfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.35
X1 XM2/vout XM2/vin VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
